`timescale 1ns / 1ps
`default_nettype none

module bmc_decoder(input wire clk, 
                   input wire [63:0] i_block,
                   output logic [63:0] o_block  
    );

    // something
    
endmodule

`default_nettype wire