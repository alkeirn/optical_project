//Clk generator module
